
module DE2_Audio_Example (
	// Inputs
	CLOCK_50,
	CLOCK_27,
	KEY,

	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	I2C_SCLK,
	SW,
	
	VGA_CLK,   														//	VGA Clock
	VGA_HS,															//	VGA H_SYNC
	VGA_VS,															//	VGA V_SYNC
	VGA_BLANK,														//	VGA BLANK
	VGA_SYNC,														//	VGA SYNC
	VGA_R,   														//	VGA Red[9:0]
	VGA_G,	 														//	VGA Green[9:0]
	VGA_B,															//	VGA Blue[9:0]
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input				CLOCK_50;
input				CLOCK_27;
input		[3:0]	KEY;
input		[6:0]	SW;
output			VGA_CLK;   				//	VGA Clock
output			VGA_HS;					//	VGA H_SYNC
output			VGA_VS;					//	VGA V_SYNC
output			VGA_BLANK;				//	VGA BLANK
output			VGA_SYNC;				//	VGA SYNC
output	[7:0]	VGA_R;   				//	VGA Red[9:0]
output	[7:0]	VGA_G;	 				//	VGA Green[9:0]
output	[7:0]	VGA_B;   				//	VGA Blue[9:0]

input				AUD_ADCDAT;

// Bidirectionals
inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;

inout				I2C_SDAT;

// Outputs
output				AUD_XCK;
output				AUD_DACDAT;

output				I2C_SCLK;

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;

wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;

// Internal Registers

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/
 
/*****************************************************************************
 *                         LAB 6 SOUNDS GO HERE                               *
 *****************************************************************************/
 
 wire [31:0] f1;
 wire [31:0] f2;
 wire [31:0] f3;
 wire [31:0] f4;
 wire [31:0] f5;
 wire [31:0] f6;
 wire [31:0] f7;
 
 
 assign f1 = 32'd96000;
 assign f2 = 32'd86000;
 assign f3 = 32'd76000;
 assign f4 = 32'd71500;
 assign f5 = 32'd64000;
 assign f6 = 32'd57000;
 assign f7 = 32'd51000;
 wire alloff;
 wire [31:0] counterout;
 
 wire c_note, d_note, e_note, f_note, g_note, a_note, b_note;
 assign c_note = SW[6];
assign d_note = SW[5];
assign e_note = SW[4];
assign f_note = SW[3];
assign g_note = SW[2];
assign a_note = SW[1];
assign b_note = SW[0];

 wire[31:0] numcyc;
	wire [31:0] thing2add;
	
wire [31:0] termc, termd, terme, termf, terg, terma, termb;
 assign termc = c_note? f1:32'b0;
 assign termd = d_note? f2:32'b0;
 assign terme = e_note? f3:32'b0;
 assign termf = f_note? f4:32'b0;
 assign termg = g_note? f5:32'b0;
 assign terma = a_note? f6:32'b0;
 assign termb = b_note? f7:32'b0;

// //use muxes, then layered add
assign numcyc = termc + termd + terme + termf + termg + terma + termb;
 
 //assign numcyc = f1*c_note + f2*d_note + f3*e_note + f4*f_note + f5*g_note + f6*a_note + f7*b_note;

 nor alloffnor(alloff, c_note, d_note, e_note, f_note, g_note, a_note, b_note);

 //assign numcyc = 32'd500000;
 
 counter audio_counter(CLOCK_50, numcyc, counterout);
 	
 assign thing2add = alloff ? 32'b0 : counterout;
 
 /*****************************************************************************
 *                         LAB 6 SOUNDS END HERE                              *
 *****************************************************************************/


assign read_audio_in			= audio_in_available & audio_out_allowed;

wire [31:0] left_in, right_in, left_out, right_out;
assign left_in = left_channel_audio_in;
assign right_in = right_channel_audio_in;


assign left_channel_audio_out	= left_out + thing2add;
assign right_channel_audio_out	= right_out + thing2add;
assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT),

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.I2C_SCLK					(I2C_SCLK),
	.I2C_SDAT					(I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0]),
	.key1							(KEY[1]),
	.key2							(KEY[2])
);

// VGA
Reset_Delay			r0	(.iCLK(CLOCK_50),.oRESET(DLY_RST)	);
VGA_Audio_PLL 		p1	(.areset(~DLY_RST),.inclk0(CLOCK_50),.c0(VGA_CTRL_CLK),.c1(AUD_CTRL_CLK),.c2(VGA_CLK)	);
vga_controller vga_ins(.iRST_n(DLY_RST),
							 .iVGA_CLK(VGA_CLK),
							 .oBLANK_n(VGA_BLANK),
							 .oHS(VGA_HS),
							 .oVS(VGA_VS),
							 .b_data(VGA_B),
							 .g_data(VGA_G),
							 .r_data(VGA_R),
							 .c(c_note),
							 .d(d_note),
							 .e(e_note),
							 .f(f_note),
							 .g(g_note),
							 .a(a_note),
							 .b(b_note));

endmodule

